module xorgate(a,b,out);
	input a,b;
	output out;
	xor(out,a,b);
endmodule
