module three_input (a,b,c,out);
	input a,b,c;
	output out;

	and(out,a,b,c);
endmodule
